module mul_matrix(clk,reset,A0,A1,A2,A3,B0,B1,B2,B3,C0,C1,C2,C3);
	input clk,reset;
	input [63:0]A0,A1,A2,A3,B0,B1,B2,B3;
	output reg [63:0]C0,C1,C2,C3;

endmodule 
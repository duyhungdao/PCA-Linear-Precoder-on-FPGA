module sq(clk,reset,x1,x2,n);
	input clk,reset;
	input [63:0] x1,x2;
	output reg [31:0]n;
endmodule
